--------------------------------------------------------------------------------
--
-- Top File for the Example Testbench (simulation)
--
--------------------------------------------------------------------------------
--
-- (c) Copyright 2009 - 2013 Advanced Micro Devices, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of Advanced Micro Devices, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- AMD, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) AMD shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or AMD had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- AMD products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of AMD products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.

--------------------------------------------------------------------------------
-- Filename: axi_bram_ctrl_0_tb.vhd
-- Description:
--  Testbench Top
--------------------------------------------------------------------------------
--
--------------------------------------------------------------------------------
-- Library Declarations
--------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

LIBRARY work;
USE work.ALL;

ENTITY axi_bram_ctrl_0_tb IS
END ENTITY;


ARCHITECTURE axi_bram_ctrl_0_tb_ARCH OF axi_bram_ctrl_0_tb IS
 SIGNAL  STATUS : STD_LOGIC_VECTOR(6 DOWNTO 0);
 SIGNAL  CLK :  STD_LOGIC := '1';
 SIGNAL  RESET : STD_LOGIC;

component axi_bram_ctrl_0_synth
PORT(
	CLK_IN     : IN  STD_LOGIC;
    RESET_IN   : IN  STD_LOGIC;
    STATUS     : OUT STD_LOGIC_VECTOR(6 DOWNTO 0) := (OTHERS => '0')   --ERROR STATUS OUT OF FPGA
    );
end component;
 
 BEGIN

  
 CLK_GEN: PROCESS BEGIN
     CLK <= NOT CLK;
     WAIT FOR 100 NS;
     CLK <= NOT CLK; 
     WAIT FOR 100 NS;
  END PROCESS;
  
  RST_GEN: PROCESS BEGIN
    RESET <= '1';
    WAIT FOR 1000 NS;
    RESET <= '0';
    WAIT;
  END PROCESS;

PROCESS BEGIN
  WAIT UNTIL STATUS(6)='1';
  IF( STATUS(5 downto 0)/="0") THEN
    ASSERT false
     REPORT "Simulation Failed"
	 SEVERITY FAILURE;
  ELSE
   ASSERT false
     REPORT "Test Completed Successfully"
	 SEVERITY FAILURE;
  END IF;
END PROCESS;	 
  
  axi_bram_ctrl_0_synth_inst: axi_bram_ctrl_0_synth
  --GENERIC MAP (
  --  C_ROM_SYNTH => 0
  --)
  PORT MAP(
           CLK_IN   => CLK,
     	   RESET_IN => RESET,
           STATUS   => STATUS
	  );

END ARCHITECTURE;
